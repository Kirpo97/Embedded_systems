`define H 4